`include "dff.v"
`include "instruction_memory.v"
`include "instructiondecoder.v"
`include ""

module CPU (
	output[1023:0] registers
);


endmodule