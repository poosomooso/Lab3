
module InstructionDecoder (
	input[31:0] instruction,
	output[5:0] opcode,
	output[4:0] rs,
	output[4:0] rt,
	output[4:0] rd,
	output[15:0] imm,
	output[25:0] addr
);



endmodule