`include "dff.v"
`include "instruction_memory.v"
`include "instructiondecoder.v"
`include "CPUcontroller.v"
`include "adder.v"
`include "alu.v"
`include "datamemory.v"
`include "signextend.v"
`include "regfile.v"


module CPU (
	output[1023:0] registers
);


endmodule